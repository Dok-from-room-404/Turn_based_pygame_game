��       ]�(KKPKe.